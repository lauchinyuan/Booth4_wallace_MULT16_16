`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Zhengzhou University
// Author: lauchinyuan
// email:lauchinyuan@yeah.net
// Create Date: 2023/04/09 16:14:57
// Module Name: tb_booth2_pp_compressor
// Description: testbench for booth2_pp_compressor Module
//////////////////////////////////////////////////////////////////////////////////


module tb_booth2_pp_compressor(

    );
    
    reg [16:0] PP1      ;
    reg [16:0] PP2      ;
    reg [16:0] PP3      ;
    reg [16:0] PP4      ;
    reg [16:0] PP5      ;
    reg [16:0] PP6      ;
    reg [16:0] PP7      ;
    reg [16:0] PP8      ;
    
    wire[30:0] PPout1   ;
    wire[28:0] PPout2   ;
    
    initial begin
        PP1 <= 17'b0_0000_0000_0000_0001;
        PP2 <= 17'b0_0000_0000_0000_0001;
        PP3 <= 17'b0_0000_0000_0000_0001;
        PP4 <= 17'b0_0000_0000_0000_0001;
        PP5 <= 17'b0_0000_0000_0000_0001;
        PP6 <= 17'b0_0000_0000_0000_0001;
        PP7 <= 17'b0_0000_0000_0000_0001;
        PP8 <= 17'b0_0000_0000_0000_0001;
    #20        
        PP1 <= 17'b0_0000_0000_0000_1001;
        PP2 <= 17'b0_0000_0000_0000_1001;
        PP3 <= 17'b0_0000_0000_0000_1001;
        PP4 <= 17'b0_0000_0000_0000_1001;
        PP5 <= 17'b0_0000_0000_0000_1001;
        PP6 <= 17'b0_0000_0000_0000_1001;
        PP7 <= 17'b0_0000_0000_0000_1001;
        PP8 <= 17'b0_0000_0000_0000_1001;   

    #20
        PP1 <= 17'b0_0000_0000_0010_1101;
        PP2 <= 17'b0_0000_0000_0010_1101;
        PP3 <= 17'b0_0000_0000_0010_1101;
        PP4 <= 17'b0_0000_0000_0010_1101;
        PP5 <= 17'b0_0000_0000_0010_1101;
        PP6 <= 17'b0_0000_0000_0010_1101;
        PP7 <= 17'b0_0000_0000_0010_1101;
        PP8 <= 17'b0_0000_0000_0010_1101;           
    end
    
    
    booth2_pp_compressor booth2_pp_compressor_inst(
        //8个部分积,这里的部分还未进行移位补零操作，
        //PP1为booth2乘数编码最低位与被乘数相乘而产生的
        //PP8为booth2乘数编码最高位与被乘数相乘而产生的
        //即PP1为做竖式乘法运算由上往下第一行
        .PP1    (PP1    ),
        .PP2    (PP2    ),  
        .PP3    (PP3    ),
        .PP4    (PP4    ),
        .PP5    (PP5    ),
        .PP6    (PP6    ),
        .PP7    (PP7    ),
        .PP8    (PP8    ),

        .PPout1 (PPout1 ),  //压缩后生成的两个部分积
        .PPout2 (PPout2 )
    );
endmodule
